-----------------------------------------------------------------------------
--
--  CPU TB constants package
--
--  This package defines constant vectors used in the CPU test bench
--
--  Revision History
--
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

package TBConstants is
    constant CLK_PERIOD : time := 20 ns;
    constant TEST_SIZE : natural := 760; -- number of clocks for test program

    type DB16Vector is array(natural range <>) of std_logic_vector(15 downto 0);
    --signal ProgABTest : DB16Vector(TEST_SIZE_AB downto 0); -- ProgAB expected output
    --signal DataABTest : DB16Vector(TEST_SIZE downto 0); -- DataAB expected output

    type DB8Vector is array(natural range <>) of std_logic_vector(7 downto 0);
	--signal DataDBWrTest : DB8Vector(TEST_SIZE downto 0); -- DataDb expected write output
    --signal DataDBRdTest : DB8Vector(TEST_SIZE downto 0); -- DataDB expected read input

    --signal DataRdTest : std_logic_vector(TEST_SIZE downto 0); -- expected data rd enable signal
    --signal DataWrTest : std_logic_vector(TEST_SIZE downto 0); -- expected data wr enable signal

    constant ProgABTest: DB16Vector(TEST_SIZE downto 0) :=(
        X"0000", X"0001", X"0002", X"0003", X"0004",
        X"0005", X"0006", X"0007", X"0008", X"0009",
        X"000A", X"000B", X"000C", X"000D", X"000E",
        X"000F", X"0010", X"0011", X"0012", X"0013",
        X"0014", X"0015", X"0016", X"0017", X"0018",
        X"0019", X"0019", X"001A", X"001B", X"001B", X"001C",
        X"001D", X"001E", X"001F", X"0020", X"0021",
        X"0022", X"0023", X"0024", X"0025", X"0026",
        X"0027", X"0027", X"0028", X"0029", X"002A", X"002B",
        X"002C", X"002D", X"002E", X"002F", X"0030", X"0030",
        X"0031", X"0032", X"0033", X"0034", X"0035",
        X"0036", X"0037", X"0038", X"0039", X"0039", X"003A",
        X"003B", X"003C", X"003D", X"003E", X"003F",
        X"0040", X"0041", X"0042", X"0043", X"0044", X"0044",
        X"0045", X"0046", X"0047", X"0048", X"0048", X"0049",
        X"004A", X"004B", X"004C", X"004D", X"004E",
        X"004F", X"0050", X"0051", X"0052", X"0053",
        X"0054", X"0055", X"0056", X"0056", X"0057", X"0058",
        X"0059", X"005A", X"005B", X"005C", X"005D",
        X"005E", X"005E", X"005F", X"0060", X"0061", X"0062",
        X"0063", X"0064", X"0065", X"0066", X"0066", X"0067",
        X"0068", X"0069", X"006A", X"006B", X"006C",
        X"006D", X"006D", X"006E", X"006F", X"0070", X"0071",
        X"0072", X"0073", X"0074", X"0075", X"0075", X"0076",
        X"0077", X"0078", X"0079", X"007A", X"007B",
        X"007C", X"007D", X"007D", X"007E", X"007F", X"0080",
        X"0081", X"0082", X"0083", X"0084", X"0085",
        X"0086", X"0086", X"0087", X"0088", X"0089", X"008A", X"008A",
        X"008B", X"008C", X"008D", X"008E", X"008E", X"008F",
        X"0090", X"0091", X"0092", X"0092", X"0093", X"0094",
        X"0095", X"0096", X"0096", X"0097", X"0098", X"0099",
        X"009A", X"009A", X"009B", X"009C", X"009D", X"009E",
        X"009F", X"009F", X"00A0", X"00A1", X"00A2", X"00A3",
        X"00A4", X"00A5", X"00A6", X"00A6", X"00A7", X"00A8",
        X"00A9", X"00AA", X"00AB", X"00AC", X"00AD",
        X"00AE", X"00AF", X"00B0", X"00B1", X"00B2",
        X"00B3", X"00B4", X"00B5", X"00B6", X"00B7", X"00B7",
        X"00B8", X"00B9", X"00BA", X"00BB", X"00BC",
        X"00BD", X"00BE", X"00BE", X"00BF", X"00C0", X"00C1",
        X"00C2", X"00C3", X"00C4", X"00C5", X"00C6",
        X"00C7", X"00C8", X"00C9", X"00CA", X"00CB",
        X"00CC", X"00CD", X"00CE", X"00CF", X"00D0",
        X"00D1", X"00D2", X"00D3", X"00D4", X"00D5",
        X"00D6", X"00D7", X"00D8", X"00D9", X"00DA",
        X"00DB", X"00DC", X"00DD", X"00DE", X"00DF",
        X"00E0", X"00E1", X"00E2", X"00E3", X"00E4",
        X"00E5", X"00E6", X"00E7", X"00E8", X"00E9",
        X"00EA", X"00EB", X"00EC", X"00ED", X"00EE",
        X"00EF", X"00F0", X"00F1", X"00F2", X"00F3",
        X"00F4", X"00F5", X"00F6", X"00F7", X"00F8",
        X"00F9", X"00FA", X"00FB", X"00FC", X"00FD",
        X"00FE", X"00FF", X"0100", X"0101", X"0102",
        X"0103", X"0104", X"0105", X"0106", X"0107",
        X"0108", X"0109", X"010A", X"010B", X"010C",
        X"010D", X"010E", X"010F", X"0110", X"0111",
        X"0112", X"0113", X"0114", X"0115", X"0116",
        X"0117", X"0118", X"0119", X"011A", X"011B",
        X"011C", X"011D", X"011E", X"011F", X"0120",
        X"0121", X"0122", X"0123", X"0124", X"0125",
        X"0126", X"0127", X"0128", X"0129", X"012A",
        X"012B", X"012C", X"012D", X"012E", X"012F",
        X"0130", X"0131", X"0132", X"0133", X"0134",
        X"0135", X"0136", X"0137", X"0138", X"0139",
        X"013A", X"013B", X"013C", X"013D", X"013E",
        X"013F", X"0140", X"0141", X"0142", X"0143",
        X"0144", X"0145", X"0146", X"0147", X"0148",
        X"0149", X"014A", X"014B", X"014C", X"014D",
        X"014E", X"014F", X"0150", X"0151", X"0152",
        X"0153", X"0154", X"0155", X"0156", X"0157",
        X"0158", X"0159", X"015A", X"015B", X"015C",
        X"015D", X"015E", X"015F", X"0160", X"0161",
        X"0162", X"0163", X"0163", X"0164", X"0165",
        X"0166", X"0167", X"0168", X"0169", X"016A",
        X"016B", X"016C", X"016D", X"016E", X"016F",
        X"0170", X"0171", X"0172", X"0173", X"0174",
        X"0175", X"0176", X"0177", X"0178",
        X"0179", X"017A", X"017B", X"017C", X"017D",
        X"017E", X"017F", X"0180", X"0180", X"0181", X"0182",
        X"0183", X"0184", X"0185", X"0185", X"0186",
        X"0187", X"0188", X"0189", X"018A", X"018B",
        X"018C", X"018D", X"018E", X"018E", X"018F",
        X"0190", X"0191", X"0192", X"0193", X"0194",
        X"0195", X"0196", X"0197", X"0197", X"0198", X"0199",
        X"0199", X"019A", X"019B", X"019C", X"019D",
        X"019E", X"019E", X"019F", X"01A0", X"01A1",
        X"01A2", X"01A3", X"01A4", X"01A5", X"01A6",
        X"01A7", X"01A7", X"01A8", X"01A9", X"01AA", X"01AB",
        X"01AB", X"01AC", X"01AD", X"01AE", X"01AF",
        X"01B0", X"01B1", X"01B2", X"01B2", X"01B3",
        X"01B4", X"01B5", X"01B6", X"01B7", X"01B7", X"01B8",
        X"01B9", X"01BA", X"01BB", X"01BB", X"01BC",
        X"01BD", X"01BE", X"01BF", X"01C0", X"01C1",
        X"01C2", X"01C2", X"01C3", X"01C4", X"01C5",
        X"01C6", X"01C7", X"01C7", X"01C8", X"01C9", X"01CA",
        X"01CB", X"01CC", X"01CC", X"01CD", X"01CE",
        X"01CF", X"01D0", X"01D1", X"01D2", X"01D3",
        X"01D4", X"01D5", X"01D5", X"01D6", X"01D7", X"01D8",
        X"01D9", X"01DA", X"01DA", X"01DB", X"01DC",
        X"01DD", X"01DE", X"01DF", X"01E0", X"01E1",
        X"01E2", X"01E3", X"01E3", X"01E4", X"01E5", X"01E5", X"01E6",
        X"01E7", X"01E8", X"01E9", X"01EA", X"01EB",
        X"01EC", X"01ED", X"01EE", X"01EF", X"01F0",
        X"01F1", X"01F2", X"01F3", X"01F4", X"01F5",
        X"01F6", X"01F7", X"01F8", X"01F9", X"01FA",
        X"01FB", X"01FC", X"01FC", X"01FD", X"01FE",
        X"01FF", X"0200", X"0201", X"0201", X"0202",
        X"0203", X"0204", X"0205", X"0206", X"0206",
        X"0207", X"0208", X"0209", X"020A", X"020B",
        X"020C", X"020D", X"020D", X"020E", X"020F",
        X"0210", X"0211", X"0212", X"0212", X"0213",
        X"0214", X"0215", X"0216", X"0217", X"0218",
        X"0219", X"0219", X"021A", X"021B", X"021C",
        X"021D", X"021E", X"021F", X"0220", X"0220",
        X"0221", X"0222", X"0223", X"0224", X"0225",
        X"0226", X"0227", X"0227", X"0228", X"0229",
        X"022A", X"022B", X"022C", X"022C", X"022D",
        X"022E", X"022F", X"0230", X"0231", X"0232",
        X"0233", X"0233", X"0234", X"0235", X"0236",
        X"0237", X"0238", X"0239", X"023A", X"023A",
        X"023B", X"023C", X"023D", X"023E", X"023F",
        X"0240", X"0241", X"0241", X"0242", X"0243",
        X"0244", X"0245", X"0246", X"0246", X"0247",
        X"0248", X"0249", X"024A", X"024B", X"024C",
        X"024D", X"024D", X"024E", X"024F", X"0250",
        X"0251", X"0252", X"0253", X"0254", X"0254",
        X"0255", X"0255", X"0256", X"0257", X"0258",
        X"0259", X"025A", X"025B", X"025C", X"025C",
        X"025D", X"025D", X"025E", X"025F", X"0260",
        X"0261", X"0262", X"0262", X"0263", X"0264", X"0264", X"0265",
        X"0266", X"0267", X"0268", X"0269", X"026A",
        X"026B", X"026C", X"026D", X"026E", X"026F",
        X"0270", X"0271", X"0272", X"0273", X"0274",
        X"0275", X"0276", X"0277", X"0278", X"0279",
        X"027A", X"027B", X"027C", X"027D", X"027E",
        X"027F", X"0280", X"0281", X"0282", X"0283",
        X"0284", X"0285", X"0286", X"0287",
        X"0289", X"028A", X"028B", X"028C", X"028D", X"028D", X"028D",--; RCALL
        X"02A1", X"02A2", X"02A3", X"02A3", X"02A3", X"02A3",
        X"028E", X"028F", X"0290", X"0291", X"0291", X"0291", -- RCALL
        X"02A1", X"02A2", X"02A3", X"02A3", X"02A3", X"02A3",
        X"0292",
        X"0293", X"0295", X"0296", X"0297",
        X"0298", X"0298", X"0298", -- ICALL
        X"02A1", X"02A2", X"02A3", X"02A3", X"02A3", X"02A3",
        X"0299", X"029A", X"029B", X"029C", X"029C", 
        X"029D", X"029D", X"029E", X"029F", X"029F", X"029F", X"029F"
    );
    constant DataABTest  : DB16Vector(TEST_SIZE downto 0) :=
    ("----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    X"FE00",            "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", X"FE00",            "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", X"FE01",            "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", X"FE02",            "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    X"FE03",            "----------------", "----------------", "----------------", "----------------",
    X"FE00",            "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    X"FF00",            "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", X"FF00",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", X"FF00",            "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", X"FF00",            "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    X"FF00",            "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", X"FF00",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", X"FF00",
    "----------------", "----------------", "----------------", "----------------", X"0070",
    "----------------", "----------------", "----------------", "----------------", X"0071",
    "----------------", "----------------", "----------------", "----------------", X"FF00",
    "----------------", "----------------", "----------------", "----------------", X"FF80",
    "----------------", "----------------", "----------------", "----------------", X"FF81",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    X"FF00",            "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", X"FF00",            "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", X"FF00",            "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", X"FF00",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", X"FF23",            "----------------", "----------------",
    "----------------", "----------------", X"FF23",            "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", X"FF23",            "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", X"FF24",            "----------------",
    X"FF24",            "----------------", "----------------", "----------------", "----------------",
    "----------------", X"FF23",            "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", X"FF45",            "----------------", "----------------",
    "----------------", X"FF45",            "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", X"FF45",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", X"FEA1",            "----------------", "----------------", "----------------",
    X"FEA1",            "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", X"FEA1",            "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    X"0076",            "----------------", "----------------", "----------------", "----------------",
    X"0076",            "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", X"FF81",            "----------------", "----------------",
    X"FF81",            "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", X"007B",            "----------------",
    "----------------", "----------------", "----------------", "----------------", X"007B",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    X"007B",            "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", X"007B",            "----------------",
    "----------------", "----------------", "----------------", "----------------", X"007A",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", X"007A",            "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    X"0069",            "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", X"0069",            "----------------",
    "----------------", "----------------", "----------------", "----------------", X"0068",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", X"0068",            "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    X"0088",            "----------------", X"0088",            "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    X"0078",            "----------------", X"0078",            "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", X"FE57",
    "----------------", "----------------", X"FE57",            "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------",
    "----------------", "----------------", "----------------", "----------------", "----------------");
    constant DataDBWrTest : DB8Vector(TEST_SIZE downto 0) :=(
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        X"00",      "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", X"01",      "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", X"02",      "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", X"34",      "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        X"1B",      "--------", "--------", "--------", "--------",
        X"0C",      "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        X"14",      "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", X"02",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", X"14",      "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", X"02",      "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        X"15",      "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", X"19",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", X"19",
        "--------", "--------", "--------", "--------", X"18",
        "--------", "--------", "--------", "--------", X"08",
        "--------", "--------", "--------", "--------", X"0A",
        "--------", "--------", "--------", "--------", X"0A",
        "--------", "--------", "--------", "--------", X"4A",
        "--------", "--------", "--------", "--------", "--------",
        X"4A",      "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", X"02",      "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", X"18",      "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", X"02",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", X"01",      "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", X"22",      "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", X"EE",      "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", X"78",      "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        X"06",      "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------",  "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", X"2B",      "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", X"58",      "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        X"12",      "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", X"44",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        X"12",      "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", X"44",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        X"73",      "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        X"73",      "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", X"99",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------", 
        "--------", "--------", "--------", "--------", "--------");

    constant DataDbRdTest : DB8Vector(TEST_SIZE downto 0) := (
        "--------", "--------", "--------", 
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", X"01",      "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", X"01",      "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        X"22",      "--------", "--------", "--------", "--------",
        "--------", X"01",      "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", X"EE",      "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", X"EE",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        X"78",      "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", X"78",      "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        X"06",      "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", X"FF",      "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        X"2B",      "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", X"58",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", X"12",      "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", X"44",      "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", X"12",      "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", X"44",      "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", X"73",      "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", X"73",      "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", X"99",      "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
        "--------", "--------", "--------", "--------", "--------",
         "--------", "--------", "--------", "--------", "--------");


    constant DataRdTest : std_logic_vector(TEST_SIZE downto 0) :=("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111011111111111101111101111111111111101111111011111111110111111101111111111101111111111111110111111111111101111111111111111111111111111011111111111110111111111111101111111111111110111111111111101111111111111110111111111111101111111110111111111011111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
    constant DataWrTest : std_logic_vector(TEST_SIZE downto 0) :=("11111111111111111111111111111101111111111110111111111011111111101111111111101111011111111111111011111111011111111011111110111111110111111110111111111011110111101111011110111101111101111111011111111111111111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111110111111111111111111011111111111111111101111111111111111110111111111111111011111111111111101111111111111111111111111011111111111011111111111110111111111111111011111111111110111111111111111011111111111110111111111111111011111111101111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

end package TBConstants;
